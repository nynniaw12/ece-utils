module ${PROJECT_NAME} (
    input  wire        clk,
    input  wire        rst_n
    // inputs + outputs
);
    // implement module
endmodule
